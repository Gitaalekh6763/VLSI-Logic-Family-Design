magic
tech scmos
timestamp 1664649723
<< nwell >>
rect 20 -10 41 22
<< polysilicon >>
rect -10 4 -8 7
rect -2 4 0 7
rect 19 4 21 7
rect 27 4 29 7
<< ndiffusion >>
rect -8 19 -2 20
rect -8 15 -7 19
rect -3 15 -2 19
rect -8 7 -2 15
rect -8 -3 -2 4
rect -8 -7 -7 -3
rect -3 -7 -2 -3
rect -8 -8 -2 -7
<< pdiffusion >>
rect 21 19 27 20
rect 21 15 22 19
rect 26 15 27 19
rect 21 7 27 15
rect 21 -3 27 4
rect 21 -7 22 -3
rect 26 -7 27 -3
rect 21 -8 27 -7
<< metal1 >>
rect -21 19 -15 20
rect 7 19 11 23
rect -21 15 -20 19
rect -16 15 -7 19
rect -3 15 22 19
rect -21 -8 -15 15
rect 34 -3 40 20
rect -3 -7 22 -3
rect 26 -7 36 -3
rect 7 -11 11 -7
rect 34 -8 40 -7
<< ntransistor >>
rect -8 4 -2 7
<< ptransistor >>
rect 21 4 27 7
<< polycontact >>
rect 0 3 4 8
rect 15 3 19 8
<< ndcontact >>
rect -7 15 -3 19
rect -7 -7 -3 -3
<< pdcontact >>
rect 22 15 26 19
rect 22 -7 26 -3
<< psubstratepcontact >>
rect -20 15 -16 19
<< nsubstratencontact >>
rect 36 -7 40 -3
<< end >>
