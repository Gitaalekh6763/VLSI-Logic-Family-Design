magic
tech scmos
timestamp 1664641249
<< nwell >>
rect -16 -3 32 12
<< polysilicon >>
rect -4 4 -1 6
rect 6 4 9 6
rect 17 4 20 6
rect -4 -26 -1 -2
rect 6 -26 9 -2
rect 17 -9 20 -2
rect 18 -13 20 -9
rect 17 -26 20 -13
rect -4 -34 -1 -32
rect 6 -34 9 -32
rect 17 -34 20 -32
<< ndiffusion >>
rect -10 -27 -4 -26
rect -10 -31 -9 -27
rect -5 -31 -4 -27
rect -10 -32 -4 -31
rect -1 -27 6 -26
rect -1 -31 1 -27
rect 5 -31 6 -27
rect -1 -32 6 -31
rect 9 -27 17 -26
rect 9 -31 11 -27
rect 15 -31 17 -27
rect 9 -32 17 -31
rect 20 -27 26 -26
rect 20 -31 21 -27
rect 25 -31 26 -27
rect 20 -32 26 -31
<< pdiffusion >>
rect -10 3 -4 4
rect -10 -1 -9 3
rect -5 -1 -4 3
rect -10 -2 -4 -1
rect -1 -2 6 4
rect 9 -2 17 4
rect 20 3 26 4
rect 20 -1 21 3
rect 25 -1 26 3
rect 20 -2 26 -1
<< metal1 >>
rect -13 8 -9 12
rect -5 8 29 12
rect -9 3 -5 8
rect 21 -18 25 -1
rect 1 -22 25 -18
rect 1 -27 5 -22
rect 21 -27 25 -22
rect -9 -36 -5 -31
rect 11 -36 15 -31
rect -13 -40 -9 -36
rect -5 -40 11 -36
rect 15 -40 29 -36
<< ntransistor >>
rect -4 -32 -1 -26
rect 6 -32 9 -26
rect 17 -32 20 -26
<< ptransistor >>
rect -4 -2 -1 4
rect 6 -2 9 4
rect 17 -2 20 4
<< polycontact >>
rect -8 -13 -4 -9
rect 2 -13 6 -9
rect 14 -13 18 -9
<< ndcontact >>
rect -9 -31 -5 -27
rect 1 -31 5 -27
rect 11 -31 15 -27
rect 21 -31 25 -27
<< pdcontact >>
rect -9 -1 -5 3
rect 21 -1 25 3
<< psubstratepcontact >>
rect -9 -40 -5 -36
rect 11 -40 15 -36
<< nsubstratencontact >>
rect -9 8 -5 12
<< end >>
