* SPICE3 file created from 3nand.ext - technology: scmos

.option scale=1u

M1000 w_n34_n9# a_3_n37# a_n14_n6# w_n34_n9# pfet w=10 l=3
+  ad=290 pd=98 as=400 ps=120
M1001 a_n14_n6# a_23_n37# a_10_n56# Gnd nfet w=10 l=3
+  ad=190 pd=58 as=170 ps=54
M1002 a_n14_n56# a_n21_n37# a_n29_n56# Gnd nfet w=10 l=3
+  ad=210 pd=62 as=120 ps=44
M1003 a_n14_n6# a_23_n37# w_n34_n9# w_n34_n9# pfet w=10 l=3
+  ad=0 pd=0 as=0 ps=0
M1004 a_10_n56# a_3_n37# a_n14_n56# Gnd nfet w=10 l=3
+  ad=0 pd=0 as=0 ps=0
M1005 a_n14_n6# a_n21_n37# w_n34_n9# w_n34_n9# pfet w=10 l=3
+  ad=0 pd=0 as=0 ps=0
C0 a_23_n37# w_n34_n9# 2.10fF
C1 a_3_n37# w_n34_n9# 2.10fF
C2 a_n21_n37# w_n34_n9# 2.10fF
C3 a_n29_n56# Gnd 18.57fF
C4 a_n14_n6# Gnd 16.36fF
C5 a_23_n37# Gnd 12.79fF
C6 a_3_n37# Gnd 12.79fF
C7 a_n21_n37# Gnd 12.79fF
