magic
tech scmos
timestamp 1664651861
<< nwell >>
rect 6 42 24 57
<< polysilicon >>
rect 28 69 31 71
rect 14 48 16 50
rect 0 34 10 38
rect 0 4 3 34
rect 14 29 16 43
rect 28 37 31 64
rect 14 22 16 24
rect 0 -3 3 -1
<< ndiffusion >>
rect -9 65 28 69
rect -13 64 28 65
rect 31 65 37 69
rect 31 64 41 65
rect 13 24 14 29
rect 16 24 17 29
rect -13 3 0 4
rect -9 -1 0 3
rect 3 3 41 4
rect 3 -1 37 3
<< pdiffusion >>
rect 13 43 14 48
rect 16 43 17 48
<< metal1 >>
rect -9 78 24 82
rect -13 69 -9 78
rect 9 52 17 56
rect 9 51 21 52
rect 9 48 13 51
rect 17 37 21 43
rect 17 33 27 37
rect 17 29 21 33
rect 9 21 13 24
rect 9 20 21 21
rect 13 16 21 20
rect 37 3 41 65
rect -13 -10 -9 -1
rect -9 -14 24 -10
<< ntransistor >>
rect 28 64 31 69
rect 14 24 16 29
rect 0 -1 3 4
<< ptransistor >>
rect 14 43 16 48
<< polycontact >>
rect 10 34 14 38
rect 27 33 31 37
<< ndcontact >>
rect -13 65 -9 69
rect 37 65 41 69
rect 9 24 13 29
rect 17 24 21 29
rect -13 -1 -9 3
rect 37 -1 41 3
<< pdcontact >>
rect 9 43 13 48
rect 17 43 21 48
<< psubstratepcontact >>
rect -13 78 -9 82
rect 9 16 13 20
rect -13 -14 -9 -10
<< nsubstratencontact >>
rect 17 52 21 56
<< end >>
