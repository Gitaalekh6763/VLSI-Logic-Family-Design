.title 3inputNOR_20bec001
.include techfile130.txt

Mp1 n1 A Vdd Vdd pmos w=260n l=130n
Mp2 n2 B n1 Vdd pmos w=260n l=130n
Mp3 Y C n2 Vdd pmos w=260n l=130n

Mn1 Y A 0 0 nmos w=130n l=130n
Mn2 Y B 0 0 nmos w=130n l=130n
Mn3 Y B 0 0 nmos w=130n l=130n

Vdd Vdd 0 1.2

VA A 0 PULSE (0 1.2 0 1n 1n 50n 100n)
VB B 0 PULSE (0 1.2 0 1n 1n 100n 200n)
VC C 0 PULSE (0 1.2 0 1n 1n 200n 400n)


.tran 0.1n 500n 0 0.1n
.control
run
plot V(A) V(B) V(C)
plot V(Y)
.endc

