* SPICE3 file created from Pass_OR.ext - technology: scmos

.option scale=1u

M1000 a_16_24# a_0_n3# w_6_42# w_6_42# pfet w=5 l=2
+  ad=25 pd=20 as=25 ps=20
M1001 a_16_24# a_0_n3# a_9_16# Gnd nfet w=5 l=2
+  ad=25 pd=20 as=25 ps=20
M1002 a_3_n1# a_16_24# a_n13_64# Gnd nfet w=5 l=3
+  ad=240 pd=116 as=205 ps=92
M1003 a_3_n1# a_0_n3# a_n13_n14# Gnd nfet w=5 l=3
+  ad=0 pd=0 as=65 ps=36
C0 a_n13_n14# Gnd 7.90fF
C1 a_9_16# Gnd 2.63fF
C2 a_0_n3# Gnd 17.82fF
C3 a_3_n1# Gnd 11.28fF
C4 a_16_24# Gnd 13.99fF
C5 a_n13_64# Gnd 7.90fF
