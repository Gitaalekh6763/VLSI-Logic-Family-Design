.title transmission_gate_20bec001
.include techfile130.txt
.include Inv.lib


**MOs d  g  s   b

Mn1 Y B A 0 nmos w=130n l=130n

Mp2 Y 1 A Vdd pmos w=260n l=130n

x1 B 1 Vdd inv

Vdd Vdd 0 1.2


VA A 0 PULSE (0 1.2 0 2n 2n 100n 200n)
VB B 0 PULSE (0 1.2 0 2n 2n 200n 300n)

Cload Y 0 70f

.tran 0.1n 500n 0 0.1n
.control
run
plot V(A) V(B)
plot V(Y)
.endc
