magic
tech scmos
timestamp 1664702285
<< nwell >>
rect -8 -5 9 7
<< polysilicon >>
rect -1 4 1 6
rect -1 -7 1 0
rect 0 -11 1 -7
rect -1 -15 1 -11
rect -1 -21 1 -19
<< ndiffusion >>
rect -3 -19 -1 -15
rect 1 -19 3 -15
<< pdiffusion >>
rect -3 0 -1 4
rect 1 0 3 4
<< metal1 >>
rect -12 8 10 11
rect -7 4 -3 8
rect 3 -15 7 0
rect -7 -24 -3 -19
rect -10 -28 -7 -24
rect -3 -28 10 -24
<< ntransistor >>
rect -1 -19 1 -15
<< ptransistor >>
rect -1 0 1 4
<< polycontact >>
rect -4 -11 0 -7
<< ndcontact >>
rect -7 -19 -3 -15
rect 3 -19 7 -15
<< pdcontact >>
rect -7 0 -3 4
rect 3 0 7 4
<< psubstratepcontact >>
rect -7 -28 -3 -24
<< labels >>
rlabel metal1 0 10 0 10 5 vdd
rlabel metal1 3 -26 3 -26 1 gnd
rlabel polycontact -3 -9 -3 -9 1 input
rlabel metal1 6 -9 6 -9 7 output
<< end >>
