.title 3inputNAND_20bec001
.include techfile130.txt


**MOs d  g  s   b

Mp1 Y A Vdd Vdd pmos w=260n l=130n
MP2 Y B Vdd vdd pmos w=260n l=130n
MP3 Y C Vdd vdd pmos w=260n l=130n

Mn1 Y A n1 0 nmos w=130n l=130n
Mn2 n1 B n2 0 nmos w=130n l=130n
Mn3 n2 C 0 0 nmos w=130n l=130n


Vdd Vdd 0 1.2

VA A 0 PULSE (0 1.2 0 1n 1n 50n 100n)
VB B 0 PULSE (0 1.2 0 1n 1n 98n 200n)
VC C 0 PULSE (0 1.2 0 1n 1n 198n 400n)


.tran 0.1n 500n 0 0.1n
.control
run
plot V(A) V(B) V(C)
plot V(Y)
.endc
