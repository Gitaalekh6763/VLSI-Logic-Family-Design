magic
tech scmos
timestamp 1664620173
<< nwell >>
rect -34 -9 54 30
<< polysilicon >>
rect -17 4 -14 6
rect 7 4 10 6
rect 27 4 30 6
rect -17 -46 -14 -6
rect 7 -46 10 -6
rect 27 -46 30 -6
rect -17 -58 -14 -56
rect 7 -58 10 -56
rect 27 -58 30 -56
<< ndiffusion >>
rect -29 -49 -17 -46
rect -29 -54 -24 -49
rect -20 -54 -17 -49
rect -29 -56 -17 -54
rect -14 -56 7 -46
rect 10 -56 27 -46
rect 30 -49 49 -46
rect 30 -54 36 -49
rect 40 -54 49 -49
rect 30 -56 49 -54
<< pdiffusion >>
rect -29 1 -17 4
rect -29 -4 -24 1
rect -20 -4 -17 1
rect -29 -6 -17 -4
rect -14 1 7 4
rect -14 -4 -4 1
rect 0 -4 7 1
rect -14 -6 7 -4
rect 10 1 27 4
rect 10 -4 17 1
rect 21 -4 27 1
rect 10 -6 27 -4
rect 30 1 49 4
rect 30 -4 36 1
rect 40 -4 49 1
rect 30 -6 49 -4
<< metal1 >>
rect -20 15 17 20
rect 21 15 51 20
rect -24 14 51 15
rect -24 1 -20 14
rect 17 1 21 14
rect -4 -25 0 -4
rect 36 -25 40 -4
rect -4 -29 40 -25
rect 36 -49 40 -29
rect -24 -66 -20 -54
rect -20 -71 51 -66
<< ntransistor >>
rect -17 -56 -14 -46
rect 7 -56 10 -46
rect 27 -56 30 -46
<< ptransistor >>
rect -17 -6 -14 4
rect 7 -6 10 4
rect 27 -6 30 4
<< polycontact >>
rect -21 -37 -17 -33
rect 3 -37 7 -33
rect 23 -37 27 -33
<< ndcontact >>
rect -24 -54 -20 -49
rect 36 -54 40 -49
<< pdcontact >>
rect -24 -4 -20 1
rect -4 -4 0 1
rect 17 -4 21 1
rect 36 -4 40 1
<< psubstratepcontact >>
rect -24 -71 -20 -66
<< nsubstratencontact >>
rect -24 15 -20 20
rect 17 15 21 20
<< end >>
