.title pass_transistor_20bec001
.include techfile130.txt
.include Inv.lib


*****************MOs d  g  s   b

Mn1 Y B A 0 nmos w=130n l=130n

Mn2 Y 1 B 0 nmos w=130n l=130n

x1 B 1 Vdd inv

Vdd Vdd 0 1.2


VA A 0 PULSE (0 1.2 0 2n 2n 100n 200n)
VB B 0 PULSE (0 1.2 0 2n 2n 198n 400n)


.tran 0.1n 500n 0 0.1n
.control
run
plot V(A) 
plot V(B)
plot V(Y)
.endc
