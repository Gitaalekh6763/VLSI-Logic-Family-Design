magic
tech scmos
timestamp 1664649509
<< nwell >>
rect -14 3 7 17
<< polysilicon >>
rect -18 30 -15 32
rect -18 -1 -15 25
rect -5 9 -2 11
rect -18 -5 -9 -1
rect -5 -12 -2 4
rect -5 -19 -2 -17
rect 8 -29 11 -5
rect 8 -36 11 -34
<< ndiffusion >>
rect -24 26 -23 30
rect -19 26 -18 30
rect -24 25 -18 26
rect -15 26 18 30
rect -15 25 22 26
rect -13 -16 -12 -12
rect -8 -16 -5 -12
rect -13 -17 -5 -16
rect -2 -16 1 -12
rect 5 -16 6 -12
rect -2 -17 6 -16
rect -24 -33 -22 -29
rect -18 -33 8 -29
rect -24 -34 8 -33
rect 11 -30 22 -29
rect 11 -34 18 -30
<< pdiffusion >>
rect -13 5 -12 9
rect -8 5 -5 9
rect -13 4 -5 5
rect -2 5 1 9
rect 5 5 6 9
rect -2 4 6 5
<< metal1 >>
rect -19 38 6 42
rect -23 37 6 38
rect -23 30 -19 37
rect -12 13 1 17
rect -12 12 5 13
rect -12 9 -8 12
rect 1 -1 5 5
rect 1 -5 8 -1
rect 1 -12 5 -5
rect -12 -21 -8 -16
rect -8 -25 6 -21
rect -22 -40 -18 -33
rect 18 -30 22 26
rect -22 -41 7 -40
rect -18 -45 7 -41
<< ntransistor >>
rect -18 25 -15 30
rect -5 -17 -2 -12
rect 8 -34 11 -29
<< ptransistor >>
rect -5 4 -2 9
<< polycontact >>
rect -9 -5 -5 -1
rect 8 -5 12 -1
<< ndcontact >>
rect -23 26 -19 30
rect 18 26 22 30
rect -12 -16 -8 -12
rect 1 -16 5 -12
rect -22 -33 -18 -29
rect 18 -34 22 -30
<< pdcontact >>
rect -12 5 -8 9
rect 1 5 5 9
<< psubstratepcontact >>
rect -23 38 -19 42
rect -12 -25 -8 -21
rect -22 -45 -18 -41
<< nsubstratencontact >>
rect 1 13 5 17
<< end >>
